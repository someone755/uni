1. vrstica: Komentar, naslov, opis ..., SPICE vse ignorira, boli njega kurac

.include ../models.inc
* komentar
* opis vezja
* tip elementa [r, c, l, m (MOS), g (bipolarni), i (tokovni vir), d (dioda)] + ime elementa [kakršenkoli tekst] + vozlišča (n1 n2 itd, + do - oz za MOS D-G-S) + parametri (1 2 ipd)
* vozlišče 0 je vedno masa

* neodvisni napetostni vir (lahko pišeš v_vin etc): vime n+ n- dc=1 sin=(offset,ampl,freq)...
* sin offset se uporabi v časovni analizi
vin 1   0   dc=0    sin=(0, 0.5, 1k)
vdd 2   0   dc=5
vss 5   0   dc=-5

* 1k...1000
* 1m...10e-3
* 1meg...10e6
* 1u...10e-6
rs  4   5   r=4371.57287525
rd  2   3   r=8k

* MOSFET: mime d g s b ime_modela par1=xx par2=yy
* bulk/substrat je ponavadi vezan na source
m1  3   1   4   4   model_nmos  w=2u    l=1u

* model NMOS tranzistorja: .model ime_modela tip_elementa [nmos, pmos, d, npn ...] p1=xx p2=yy
.model  model_nmos   nmos    vto=1.4    kp=0.25m
* parameter je vedno kp, za nmos ALI za pmos

* ukazi: cd, echo, op, setplot, destroy, display, print, let, dc, plot, max, min, tran
.control
destroy all
echo ###########################
echo ----------- OP1 -----------
op
let vgsq = v(1,4)
let vdsq = v(3,4)
let idq=-vdd#branch
* ali let idq=-i(vdd) -- tok skozi element

* napetostni vir z dc=0 je kratek stik, ampak lahko izmerimo tok i skozenj

print vgsq vdsq idq v(3)


echo ----------- DC1 -----------
* DC analiza: dc    ime_parametra   start   stop    korak
dc  vin -10 10  0.01

let id = -i(vdd)
let vds = v(3,4)

* plot y_os vs x_os title 'text' xlabel 'text' ylabel 'text'
* default x_os je sweep (poglej v 'display')
plot id vs vds xlabel 'vds [V]' ylabel 'id [A]'
plot v(3)

echo ---------- TRAN1 ----------
* Time-domain analysis
* čas. analiza: tran začetni_korak čas_analize začetek_shranjevanja
* tran dt tstop
tran    1u 10m

let vin=v(1)
let vout=v(3)

let vin_pp = max(vin) - min(vin)
let vout_pp = max(vout) - min(vout)
let av_abs = vout_pp/vin_pp
print av_abs * -1

plot vin vout ylabel 'r: vin[V], g:vout[V]' xlabel 't'
* setplot
* display - pokaže kaj je zračunal v zadnji analizi
* plot v(1) v(3)

* fourier: fourier  f0  signal
fourier 1k  vout

.endc

.end
