Vaja 3: MOSFET kaskodni ojačevalnik

vin	1	0	dc=0	sin(0,	0.0402,	5k)
vp	2	0	dc=5
vn 	5	0	dc=-5
* preverjanje IDQ z napetostnim virom dc=0
vcurr	7	8	dc=0
* preverjanje I_izhodni z napetostnim virom dc=0
vcurr_out	6	10	dc=0

r1	2	3	r=40483.7
r2	3	4	r=31627.9
r3	4	5	r=54400

rd	2	6	r=5k
rs	9	5	r=5k

c1	1	4	c=100u
c2	3	0	c=100u
c3	9	0	c=100u

m1	8	4	9	9	model_nmos w=1u 	l=1u
m2	6	3	7	7	model_nmos w=1u 	l=1u

.model model_nmos	nmos 	vto=0.8	kp=1m	lambda=1e-4

.control
destroy all

echo ------- OP1 -------
op
let vdsq2 = v(6,7)
let vgsq2 = v(3,7)

let vdsq1 = v(8,9)
let vgsq1 = v(4,9)

let vg1 = v(4)

let idq = vcurr#branch

print vgsq1 vgsq2 vdsq1 vdsq2 idq vg1

echo
echo ------ TRAN1 ------
tran 1u 1m

let vin = v(1)
let vout = v(6)

plot vin vout
let vin_pp = max(vin) - min(vin)
let vout_pp = max(vout) - min (vout)
let av_abs = vout_pp/vin_pp

print -av_abs

echo
echo ------ FREQ1 ------
fourier	5k	vout

echo
echo - INPUT IMPEDANCE -
let iin_pp = max(vin#branch) - min(vin#branch)
let uin_pp = max(vin) - min(vin)
let rin = uin_pp/iin_pp
print rin

.endc
.end